module Vivid.Scene.Camera

class GameCamera : GameScript

    func GameCamera()

    end 

end 