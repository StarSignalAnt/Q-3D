module Vivid.Game

class #NAME#

    func #NAME#()

    end

    func Update(float delta)

    end 

end 
