module Vivid.Game

class GameScript

    Node node;
    Input input;

    func GameScript()

        node = new Node();
        input = new Input();
        Debug("Game Script!");

    end 

  

end     